



//=================================================
// Main for tb
//=================================================
initial begin:INIT_ROM
    rom_data[0] = 256'd8373472657281772018911143333458316925033721577737104126053548254730873694134;
    rom_data[1] = 256'd7077606502272555644217196429706292779513133638075460940993818609581453840285;
    rom_data[2] = 256'd7114136467605830164386765627892048130214786415103409736546034808857167887507;
    rom_data[3] = 256'd4242306337368971763956605508238427748907152257205517154330783395676974510220;
    rom_data[4] = 256'd231497681911891134178994672965761884324664899027051010815610961774572168814;
    rom_data[5] = 256'd2519209966448930701014592276617105726045457045240388104133533414463254742751;
    rom_data[6] = 256'd6039381731594839481832183287375266550233822026911004676411544779179579562275;
    rom_data[7] = 256'd4690871450214802552634031731879642285788537203250678175927475536301984849125;
    rom_data[8] = 256'd7975009210824794677566260793836397350585861665209360099794990688301299962401;
    rom_data[9] = 256'd467620823670762988783146281724334162048150830781734579065395991105808182671;
    rom_data[10] = 256'd6107215824437711227292024781347992340585139264873923923588781987862688777840;
    rom_data[11] = 256'd5365539456217618198023417874642539899492225210021410152464686338449142766690;
    rom_data[12] = 256'd3325620720463859217255678259367663152094527211798586531628394533097127461168;
    rom_data[13] = 256'd4557410224557902980968787359427463221169015279818015765337231467258424517896;
    rom_data[14] = 256'd5942418366679351008921318488178368716010252409631424771254318350414889877990;
    rom_data[15] = 256'd2783850377373548791149416652758502964325697351893678513423050070505381001072;
    rom_data[16] = 256'd328024486901120694958175617147608978617507250200945349318384805620294159463;
    rom_data[17] = 256'd8197005208467186304575826513426424464378461765442898631363620698768737903366;
    rom_data[18] = 256'd5372281487070429983030750203387831824028937311011922850553868166709400313814;
    rom_data[19] = 256'd2606947917178271102153189518251525217685411797315460077954840610637138564973;
    rom_data[20] = 256'd3026075928655997184998462090118109524134371799196606845392710202991007379636;
    rom_data[21] = 256'd7554044695149057488166319800012513140304227924998636579758602585243216296444;
    rom_data[22] = 256'd1366243870743353208258125244342968546165415649396178220925670514214854489559;
    rom_data[23] = 256'd4997109254876689809032723042751339706315204041169791759879685098173744064999;
    rom_data[24] = 256'd424349897640303839737150584238876656973747313339179409974220601118948844933;
    rom_data[25] = 256'd1392368661687672140736515737058342795560990007760791982514243765005727830480;
    rom_data[26] = 256'd4695395786108323772524156838850626329552681302709486893249983465561221665847;
    rom_data[27] = 256'd8144810879780247726054624022948720944256855235141394716513811699310511305495;
    rom_data[28] = 256'd2288833553330634569603301341875273410674857365188490713627003364280329224085;
    rom_data[29] = 256'd5764412680380118956796127884937678993110359157540092248573201494945797828714;
    rom_data[30] = 256'd5315628833519211749819786394473370143014847532141022294747025020483061503504;
    rom_data[31] = 256'd2812552823302879012035658606070183634911359839168061409582453158348139842894;
    rom_data[32] = 256'd4689781612658861830718587139225427027672044485884334513034660528191039868271;
    rom_data[33] = 256'd3689534145322975739667156060455335418048340885547481722298563155371571699225;
    rom_data[34] = 256'd7725887051664955468679986393530293421926645356214259363050711732886927038154;
    rom_data[35] = 256'd3946289232403687999941280644147403847117686951759674818057486446459205438811;
    rom_data[36] = 256'd5579784820146992624646930169972337511846200153900265026403014092733541670449;
    rom_data[37] = 256'd3699682967984877782651937473939865099953763193116412734750712861668302978953;
    rom_data[38] = 256'd5172806624402906048472383367905622939253798645831621441907443721731869825048;
    rom_data[39] = 256'd7507592971378093139413072722528931995474572691977348966310144477230019826348;
    rom_data[40] = 256'd245134702730808611856421032763291201650792984808587875251338056482221016740;
    rom_data[41] = 256'd6465194219743152961334836997164554609332752385943418448022734533549155795953;
    rom_data[42] = 256'd7162429293317993669842002635616889614808303192269165618542497657118713317397;
    rom_data[43] = 256'd3331498932099424038563638195884719018116040974483729872803380454138162302849;
    rom_data[44] = 256'd6282051498390224539895546021249470851417154232196182350507190107264091281489;
    rom_data[45] = 256'd6813614447854539501990287843726853845514363910307187928751351556038669339809;
    rom_data[46] = 256'd5903907811897009872569783482940876163884870493678917782402512767435761648614;
    rom_data[47] = 256'd6862044436047110472825051773692380431642054209480723254226076711098277692607;
    rom_data[48] = 256'd3157305792208799014342159403356446589767965270948137452277654410355539325615;
    rom_data[49] = 256'd8212417329780623740409146145961247663469924470978880191286969542933205651012;
    rom_data[50] = 256'd5418044532993552291074858747209209318708205188166481050413166077254899985205;
    rom_data[51] = 256'd2793919512847324028906394140097535576647992698377015791548161020439271240147;
    rom_data[52] = 256'd4729622605399328650372774795544529985626493278974787246598578188728434064424;
    rom_data[53] = 256'd8377272167102186543054395652762896868516679540447826038119312832908613185254;
    rom_data[54] = 256'd1720086019607897279769638140398961561660541550467184869480709335530695533565;
    rom_data[55] = 256'd6889201701715011230093237733165279201552540041547450035271952680898736274814;
    rom_data[56] = 256'd3360301915849272161769760848002967324400322516485937307304066261469762384714;
    rom_data[57] = 256'd257305868634842875615041361830240252729191592111857522061299453353994298464;
    rom_data[58] = 256'd2997740921023779705085531090816465712895533337160786998297964010747270129913;
    rom_data[59] = 256'd153757039166444162121572512371540332299736024488228473841844465330537371715;
    rom_data[60] = 256'd48330922093538503367073388766111442406990470700873498744048821883979391792;
    rom_data[61] = 256'd3125237263893215904492512646644502899918512636369452419842214659044816475650;
    rom_data[62] = 256'd1438077745239161803715139624582066309439624948297296918545955597763320431251;
    rom_data[63] = 256'd2893324476580958220512544739216086603177004936502518340923742459413793141866;
    rom_data[64] = 256'd5668022560815707471346210357486645758873687610926719876060611915518553245070;
    rom_data[65] = 256'd2890303749660010388456593992383638639799689993495962333269169226586288946560;
    rom_data[66] = 256'd6985777019057367388925625543013425340409544870300922550978302633310479256135;
    rom_data[67] = 256'd7703831121808264771824986893499183209930502129514484562644446040426640282901;
    rom_data[68] = 256'd4275739633570171454861271688346850183849412075611304650787025237412838043272;
    rom_data[69] = 256'd1057531793335316837904295944464123732476231748240232521385227397145276753955;
    rom_data[70] = 256'd7900524496030609176318108850381374477290295981618729557380358155153561794470;
    rom_data[71] = 256'd3945351296563897506743333586190573845009416725772711243115456724413694916596;
    rom_data[72] = 256'd2141258122740212607832504011750741308071657807837895806677453167680975750603;
    rom_data[73] = 256'd591418045400760767074750787335610461670102645464781336133818048829705991091;
    rom_data[74] = 256'd5270357908433524870835701350428651770135695076327423190385074984755541469601;
    rom_data[75] = 256'd3199329410674350949662219611971363510887833464985389664699747787364826147172;
    rom_data[76] = 256'd2142669515282495747573665649182684987465738337145268990586108456118282436130;
    rom_data[77] = 256'd7705861193047179589219928696944765740688728932822735735844659092432714050498;
    rom_data[78] = 256'd4065523259541523209812128784885096957309095261079677627654826928456184811469;
    rom_data[79] = 256'd7957161268925551669358142424760511793305279760605271573010011426519013251855;
    rom_data[80] = 256'd4218140435052384771717575495961105624815706011550786329850432777261151191688;
    rom_data[81] = 256'd4840577668689279979598991558708315152548819680861494981814870214093439251617;
    rom_data[82] = 256'd6378340912455226800923521210856591952989675708848505399009200939400500737242;
    rom_data[83] = 256'd7023288836843702057298730433493858395997646534702484903144270024343232564331;
    rom_data[84] = 256'd1578820218489100815636262291641385545236341295785424626901679803901388305941;
    rom_data[85] = 256'd1567800108808253310626099447301436492994619508946411805598756878398291363117;
    rom_data[86] = 256'd2151734034940868241820000095278287899344438590418544639934490920928523395969;
    rom_data[87] = 256'd8411547382793484865074667901576255416071463179072892440732899472999046063099;
    rom_data[88] = 256'd3897192943195137482630118206349048052371533787235756220898283367759544509451;
    rom_data[89] = 256'd4957609844880988207568496253129906536580209878898248702983040607721960833431;
    rom_data[90] = 256'd1792799086573295671856704501668717172927784565556129774941459946445725125648;
    rom_data[91] = 256'd391810143215968393343828566400337584863803262665241114578787306656609196564;
    rom_data[92] = 256'd608775887523418242345898808567808596308508167354314274264323701125617011977;
    rom_data[93] = 256'd1764566075909582564316017125839334776682549089564593806545761989686334857625;
    rom_data[94] = 256'd1740775745857789223508916790664481194837782792876359783912243542018621110161;
    rom_data[95] = 256'd7912572937193886952699577425102737753579778402438476027626150530907806356615;
    rom_data[96] = 256'd3704872392311763585336177554837998539081315019618456242102333484022912807319;
    rom_data[97] = 256'd8402346693307336048694008664497015103626743700452894277236439838778131383612;
    rom_data[98] = 256'd7300348668782676956861213748488086204812414066580579682612456732180040403681;
    rom_data[99] = 256'd3462508604217227799880787078817121185613687048547043365467643451111762290437;
    rom_data[100] = 256'd4924658466610466496858396199653680606259481438444767365731834592767292380687;
    rom_data[101] = 256'd3042270273118384162682923856075540061809821163454768737682565903459292482049;
    rom_data[102] = 256'd5893165840519852158574086435438793419299529932629124229543186003828927985782;
    rom_data[103] = 256'd6207054488551387381207998415311196576842426645742482130013600028020893859801;
    rom_data[104] = 256'd4084187408678960277972350057794732238592768938562746451368356055556161711572;
    rom_data[105] = 256'd2859262363561906608311935440467932616284054493021877033117206957756241601088;
    rom_data[106] = 256'd3893097338298960378294412938640885774983770300331564614824386510926062391793;
    rom_data[107] = 256'd1629918156339470079737370175165340212398299264249646088828615758793353623247;
    rom_data[108] = 256'd1063846543378727076227610240694088876187064801378696460327862866571236024337;
    rom_data[109] = 256'd4690795036151477377422852585907129739232979379919730811301371129679125794935;
    rom_data[110] = 256'd5484569803959182588242765469608234636947834418544853369836723130527616933915;
    rom_data[111] = 256'd5520436455190686128316520374622382595982341089923365509990418823683134388711;
    rom_data[112] = 256'd7183694964249559039514553830595092487925710083298946148948449795387697569979;
    rom_data[113] = 256'd6238926434346313818359711273546319521783356418260834172711777786879398669587;
    rom_data[114] = 256'd5786191127154750903951729281367309657375886226506629629533609983720108872308;
    rom_data[115] = 256'd6918787362911162389603288270671352938456461614784584983691156381344138264730;
    rom_data[116] = 256'd4213334538681476500073322967009096853628850440431678438463496991915364647908;
    rom_data[117] = 256'd7682146375945287813431141161467080846433474287583722732393525331420980771572;
    rom_data[118] = 256'd7793341030119038627864777610284226988303618642758151649744897628206172882671;
    rom_data[119] = 256'd4379966993945925230070795483854641949318351848004236292715200553859640388605;
    rom_data[120] = 256'd4270497961777455662303735356522368200818947943945388945647374653984222296613;
    rom_data[121] = 256'd7905376038939465331349267244972492532156645071079150915867657851875634180578;
    rom_data[122] = 256'd4258089265303226495954002121419092553650549362885040057035240789194877950609;
    rom_data[123] = 256'd4508908533977769458527940766359918758512953590702270080064549950812452446332;
    rom_data[124] = 256'd213513894764764919418617042602041241975091434278342765409671444806256485227;
    rom_data[125] = 256'd7972775708699191793783629420185304001001479343330193920517094140212651080056;
    rom_data[126] = 256'd5781546459391152824522043249423532371962371676315090884479078868371754154833;
    rom_data[127] = 256'd235310776455809857314800037131144696261018915686867407678697043723786760521;
end



integer i = 0;


/*
initial
begin:UL_REQ_GEN
 @(posedge i_rst_n)
    repeat(3)
  begin
    #6us;
    @(posedge i_clk)
    ul_req = 1'b1;
    @(posedge i_clk)
    ul_req = 1'b0;

  end // end repeat
end
*/









// bfm inst

soc_cfg_send_if u_soc_if(i_clk, i_rst_n);
soc_cfg_sender sender;


assign o_last_no_rom = SVT_top.u_ped64_top_wrapper.o_last_ped64;

always@(o_last_no_rom)
  broadcast_addr = 32'h0001_0000;


  initial begin:SOC_CFG_SENDER_GEN
    broadcast_addr = 32'h0001_0000;
    `ifdef PREDICTABLE_DATA 
    //=================================================
    // Generate predictable data pattern
    // Each 32-bit word increases by +1
    // Total 8 * 256 bits = 64 * 32-bit words
    //=================================================
    bit [31:0] base = 32'h0000_0000;
    for (int blk = 0; blk < 8; blk++) begin
      for (int w = 0; w < 8; w++) begin
        soc_data_arr[blk][w*32 +: 32] = base;
        base += 1;
      end
    end
    `endif // end of PREDICTABLE_DATA

    sender = new(u_soc_if);
    while(1)
    begin
      // req
      wait(soc_req)
      
      `ifndef PREDICTABLE_DATA
      
      soc_data_arr[0]  = swap_32bit_blocks(rom_data[broadcast_addr[7:0]*2]);
      soc_data_arr[1]  = swap_32bit_blocks(rom_data[broadcast_addr[7:0]*2+1]);
      $display("[%0t] INFO: broadcast_addr = %0h ,arr_x = %0h,arr_y = %0h", $time, broadcast_addr,soc_data_arr[0],soc_data_arr[1] );
      `endif
      sender.send(broadcast_addr, soc_data_arr);
      broadcast_addr = broadcast_addr + 1'b1;
    end
  end



